module RAM_512x16_3 (
    input [8:0] ram_addr,
    input [15:0] ram_wdata,
    output [15:0] ram_rdata,
    input ce,
    input clk,
    input we,
    input re);

    wire [15:0] ram_rdata0;
    wire [15:0] ram_rdata1;

    assign ram_rdata = ram_addr[8] ? ram_rdata1 : ram_rdata0;

    SB_RAM40_4K RAM_inst0(
        .RDATA(ram_rdata0),
        .RADDR({3'b000,ram_addr[7:0]}),
        .RCLK(clk),
        .RCLKE(re&ce),
        .RE(re&ce),
        .WDATA(ram_wdata),
        .WADDR({3'b000,ram_addr[7:0]}),
        .WCLK(clk),
        .WCLKE(we&ce),
        .WE(we&ce),
        .MASK(16'h0000));
    defparam RAM_inst0.READ_MODE =0;
    defparam RAM_inst0.WRITE_MODE =0;

    SB_RAM40_4K RAM_inst1(
        .RDATA(ram_rdata1),
        .RADDR({3'b000,ram_addr[7:0]}),
        .RCLK(clk),
        .RCLKE(re&ce),
        .RE(re&ce),
        .WDATA(ram_wdata),
        .WADDR({3'b000,ram_addr[7:0]}),
        .WCLK(clk),
        .WCLKE(we&ce),
        .WE(we&ce),
        .MASK(16'h0000));
    defparam RAM_inst0.READ_MODE =0;
    defparam RAM_inst0.WRITE_MODE =0;

    /*strings*/
    defparam RAM_inst0.INIT_0 = 256'h57F2_5C64_6124_6612_6B0A_6FE8_748B_78D4_7CAB_7FFD_82C0_84F2_8698_87C2_8883_88F6;
    defparam RAM_inst0.INIT_1 = 256'h3C59_3F53_41A0_434D_4473_4530_45A7_4600_4663_46F6_47DA_492C_4B02_4D68_5062_53EA;
    defparam RAM_inst0.INIT_2 = 256'h027F_00AB_0000_0085_0236_0500_08C5_0D5F_129E_184F_1E3C_2430_29F7_2F66_3457_38AE;
    defparam RAM_inst0.INIT_3 = 256'h3A1F_3AD2_3AD8_3A14_3874_35F1_3291_2E67_2991_2439_1E90_18CF_1330_0DF0_0948_0569;
    defparam RAM_inst0.INIT_4 = 256'h31B4_313C_3090_2FCC_2F0C_2E70_2E12_2E0A_2E65_2F2B_3056_31D7_3396_3572_3744_38E1;
    defparam RAM_inst0.INIT_5 = 256'h3AB9_3645_3283_2F8D_2D6C_2C1E_2B92_2BAA_2C45_2D37_2E56_2F7A_307E_3146_31C0_31E4;
    defparam RAM_inst0.INIT_6 = 256'h5588_5807_5AB1_5D37_5F4F_60B9_6143_60CB_5F43_5CAF_5926_54CE_4FDA_4A85_450F_3FB7;
    defparam RAM_inst0.INIT_7 = 256'h8855_87E1_8583_8182_7C3A_7612_6F77_68D5_6292_5D04_5870_5507_52E0_51FB_5240_5383;
    defparam RAM_inst0.INIT_8 = 256'h0347_04F5_08EF_0F25_176A_2178_2CEF_395F_464A_532D_5F83_6AD4_74B2_7CC5_82CF_86AB;
    defparam RAM_inst0.INIT_9 = 256'h4812_49C8_4A3F_494E_46E2_42FF_3DBD_374D_2FF6_280D_1FF9_1825_1104_0B01_0681_03D8;
    defparam RAM_inst0.INIT_A = 256'h51E8_49DB_4281_3C17_36CF_32D0_302F_2EF5_2F14_3071_32DD_361D_39E8_3DEE_41DA_4556;
    defparam RAM_inst0.INIT_B = 256'h8C08_8EAA_90DA_926E_933C_931D_91F3_8FAA_8C36_879A_81E5_7B35_73B1_6B8D_6308_5A64;
    defparam RAM_inst0.INIT_C = 256'h5F6F_6392_673B_6A70_6D3E_6FBB_71FF_7425_7648_787F_7ADC_7D69_8028_8313_8619_8921;
    defparam RAM_inst0.INIT_D = 256'h2D4E_2B65_2A38_29E5_2A7D_2C08_2E81_31D8_35F1_3AAB_3FDB_4556_4AEF_5079_55D0_5AD4;
    defparam RAM_inst0.INIT_E = 256'h4C03_4AC0_49DF_4938_489E_47EA_46F8_45AC_43F6_41D0_3F3F_3C54_392D_35ED_32BF_2FD0;
    defparam RAM_inst0.INIT_F = 256'h9720_94CC_9159_8CE3_8792_8196_7B29_7484_6DE1_677A_617F_5C18_5763_536F_5041_4DCE;

    defparam RAM_inst1.INIT_0 = 256'h6CCB_6D3D_6E91_70C1_73BB_7764_7B97_8025_84DC_8982_8DDE_91B5_94D5_970E_983C_9846;
    defparam RAM_inst1.INIT_1 = 256'h9A1B_97F9_958F_92D7_8FD0_8C7F_88EE_852B_814E_7D70_79B0_762E_730E_7071_6E76_6D37;
    defparam RAM_inst1.INIT_2 = 256'hB2E6_B1AE_B041_AEB0_AD08_AB56_A9A7_A803_A66F_A4ED_A37B_A212_A0AA_9F38_9DAE_9BFE;
    defparam RAM_inst1.INIT_3 = 256'hA5E8_A696_A79D_A8F1_AA7E_AC2E_ADEA_AF9C_B12C_B288_B39E_B461_B4CA_B4D6_B484_B3DC;
    defparam RAM_inst1.INIT_4 = 256'hB28E_B334_B370_B33F_B2A4_B1AA_B060_AEDB_AD32_AB80_A9DF_A866_A72E_A647_A5C0_A5A0;
    defparam RAM_inst1.INIT_5 = 256'hB096_AD84_AAEB_A8DA_A75C_A673_A61F_A655_A708_A824_A990_AB32_ACEC_AE9F_B031_B188;
    defparam RAM_inst1.INIT_6 = 256'hE462_E2DC_E114_DF04_DCA7_D9FA_D6FE_D3B4_D023_CC53_C852_C431_C003_BBDE_B7DA_B410;
    defparam RAM_inst1.INIT_7 = 256'hDEFC_E14E_E353_E506_E66A_E781_E84F_E8D9_E926_E939_E919_E8C8_E848_E79A_E6BC_E5AB;
    defparam RAM_inst1.INIT_8 = 256'hBCA8_BBCA_BB92_BBFE_BD06_BE9F_C0B8_C33D_C61A_C938_CC7E_CFD7_D32D_D66B_D980_DC5F;
    defparam RAM_inst1.INIT_9 = 256'hEB12_EA1E_E88E_E66B_E3C2_E0A2_DD21_D957_D560_D158_CD5F_C992_C60D_C2EC_C044_BE29;
    defparam RAM_inst1.INIT_A = 256'hBE11_C243_C683_CAC4_CEFA_D318_D712_DAD9_DE60_E197_E471_E6E0_E8D4_EA44_EB22_EB69;
    defparam RAM_inst1.INIT_B = 256'hA05D_9FB3_9F45_9F20_9F50_9FDE_A0D0_A22B_A3EE_A618_A8A4_AB8C_AEC6_B248_B608_B9F9;
    defparam RAM_inst1.INIT_C = 256'hADC7_ACB1_ABCA_AB07_AA5E_A9C2_A927_A885_A7D3_A70C_A62E_A53C_A43A_A331_A22B_A135;
    defparam RAM_inst1.INIT_D = 256'hD301_D133_CF15_CCB4_CA1B_C75A_C480_C19A_BEB9_BBEC_B940_B6C1_B478_B26B_B0A0_AF14;
    defparam RAM_inst1.INIT_E = 256'hB524_B9F4_BE90_C2E4_C6E0_CA77_CD9E_D04E_D282_D437_D56E_D627_D667_D630_D588_D476;
    defparam RAM_inst1.INIT_F = 256'h8939_896C_89B1_8A26_8AE8_8C0E_8DA9_8FC7_926A_9591_9935_9D46_A1B3_A665_AB44_B037;



endmodule

